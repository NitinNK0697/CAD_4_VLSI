package int8_mac_pipe;

    interface Ifc_int8;
        method Action       put(Bit#(8) a, Bit#(8) b, Bit#(32) c);
        method Bit#(32)     get();
    endinterface

    module mk_Test(Empty);
        Reg#(int)           count <- mkReg(1);
        Reg#(Int#(8))       rg_a  <- mkReg(100);        
        Reg#(Int#(8))       rg_b  <- mkReg(100);
        Reg#(Int#(32))      rg_c  <- mkReg(500);

        Ifc_int8 obj_mac <- mk_int8_mac;

        rule inp(count==1);
            obj_mac.put(pack(rg_a),pack(rg_b),pack(rg_c));
            count <= count+1;
        endrule

        rule stall(count < 11 && count>1);
            count <= count+1;
        endrule

        rule res;
            Int#(32) rg_m = unpack(obj_mac.get());
          //  $display("Inputs: %d, %d, %d", rg_a, rg_b, rg_c);
            $display("%d  INT8 MAC O/P: %d",count, rg_m);
        endrule

        rule stop(count==11);
            $finish(0);
        endrule

    endmodule

    
// //Test Bench
//   module mk_Tb(Empty);
//     Reg#(Bit#(16)) rg_a  <- mkReg(?);        
//     Reg#(Bit#(16)) rg_b  <- mkReg(?);
//     Reg#(Bit#(32)) rg_c  <- mkReg(?);
//     Reg#(Bit#(32)) rg_mac  <- mkReg(?);
//     Reg#(Bit#(1))  rg_r  <- mkReg(1'b1);
//     Reg#(Int#(32))  count  <- mkReg(0);
//     Reg#(Int#(32))  failed_cases  <- mkReg(0);

//     Reg#(Bit#(16)) rg_af <- mkReg(?);        
//     Reg#(Bit#(16)) rg_bf <- mkReg(?); //unpack({1'b1, 8'd0, 23'd0})
//     Reg#(Bit#(32)) rg_cf <- mkReg(?);
//     Reg#(Bit#(32)) rg_macf  <- mkReg(?);

//     Reg#(Bit#(16)) as1 <- mkReg(?);
//     Reg#(Bit#(16)) bs1 <- mkReg(?);
//     Reg#(Bit#(32)) cs1 <- mkReg(?);
//     Reg#(Bit#(32)) cs2 <- mkReg(?);
//     Reg#(Bit#(32)) cs3 <- mkReg(?);
//     Reg#(Bit#(32)) cs4 <- mkReg(?);
//     Reg#(Bit#(32)) cs5 <- mkReg(?);
//     Reg#(Bit#(32)) cs6 <- mkReg(?);
//     Reg#(Bit#(32)) cs7 <- mkReg(?);
//     Reg#(Bit#(32)) cs8 <- mkReg(?);
//     Reg#(Bit#(32)) cs9 <- mkReg(?); 
//     Reg#(Bit#(16)) as2 <- mkReg(?);
//     Reg#(Bit#(16)) bs2 <- mkReg(?);
//     Reg#(Bit#(16)) as3 <- mkReg(?);
//     Reg#(Bit#(16)) bs3 <- mkReg(?);
//     Reg#(Bit#(16)) as4 <- mkReg(?);
//     Reg#(Bit#(16)) bs4 <- mkReg(?);
//     Reg#(Bit#(16)) as5 <- mkReg(?);
//     Reg#(Bit#(16)) bs5 <- mkReg(?);
//     Reg#(Bit#(16)) as6 <- mkReg(?);
//     Reg#(Bit#(16)) bs6 <- mkReg(?);
//     Reg#(Bit#(16)) as7 <- mkReg(?);
//     Reg#(Bit#(16)) bs7 <- mkReg(?);
//     Reg#(Bit#(16)) as8 <- mkReg(?);
//     Reg#(Bit#(16)) bs8 <- mkReg(?);
//     Reg#(Bit#(16)) as9 <- mkReg(?);
//     Reg#(Bit#(16)) bs9 <- mkReg(?); 
//     Reg#(Bit#(16)) as10 <- mkReg(?);
//     Reg#(Bit#(16)) bs10 <- mkReg(?);
//     Reg#(Bit#(32)) cs10 <- mkReg(?); 
//     Reg#(Bit#(16)) as11 <- mkReg(?);
//     Reg#(Bit#(16)) bs11 <- mkReg(?);
//     Reg#(Bit#(32)) cs11 <- mkReg(?);  
//     Reg#(Bit#(16)) as12 <- mkReg(?);
//     Reg#(Bit#(16)) bs12 <- mkReg(?);
//     Reg#(Bit#(32)) cs12 <- mkReg(?);

//     Reg#(Bit#(32)) macs1 <- mkReg(?);
//     Reg#(Bit#(32)) macs2 <- mkReg(?);
//     Reg#(Bit#(32)) macs3 <- mkReg(?);
//     Reg#(Bit#(32)) macs4 <- mkReg(?);
//     Reg#(Bit#(32)) macs5 <- mkReg(?);
//     Reg#(Bit#(32)) macs6 <- mkReg(?);
//     Reg#(Bit#(32)) macs7 <- mkReg(?);
//     Reg#(Bit#(32)) macs8 <- mkReg(?);
//     Reg#(Bit#(32)) macs9 <- mkReg(?);
//     Reg#(Bit#(32)) macs10 <- mkReg(?);
//     Reg#(Bit#(32)) macs11 <- mkReg(?);
//     Reg#(Bit#(32)) macs12 <- mkReg(?);
    
//     Ifc_int8 mac <- mk_int8_mac;  
//     Ifc_inp obj_inp <- mk_inp_read;        

//     rule inp;
//          obj_inp.put_r(1'b1);
//          Bit#(8) a = obj_inp.get_a();
//          Bit#(8) b = obj_inp.get_b();
//          Bit#(32) c = obj_inp.get_c();
//          Bit#(32) mac1 = obj_inp.get_mac();
//          mac.put(a,b,c);
//          rg_af <= unpack({8'd0,a});
//          rg_bf <= unpack({8'd0,b});
//          rg_cf <= unpack(c);
//          rg_macf <= unpack(mac1);
//          count <= count+1;
//     endrule


//     rule pipe;
//         //$display("Count: %d --A: %b", count, pack(rg_af));
//         as1 <= rg_af;
//         bs1 <= rg_bf;
//         cs1 <= rg_cf;
//         macs1 <= rg_macf;
//         as2 <= as1;
//         bs2 <= bs1;
//         cs2 <= cs1;
//         macs2 <= macs1;
//         as3 <= as2;
//         bs3 <= bs2;
//         cs3 <= cs2;
//         macs3 <= macs2;
//         as4 <= as3;
//         bs4 <= bs3;
//         cs4 <= cs3;
//         macs4 <= macs3;
//         as5 <= as4;
//         bs5 <= bs4;
//         cs5 <= cs4;
//         macs5 <= macs4;
//         as6 <= as5;
//         bs6 <= bs5;
//         cs6 <= cs5;
//         macs6 <= macs5;
//         as7 <= as6;
//         bs7 <= bs6;
//         cs7 <= cs6;
//         macs7 <= macs6;
//         as8 <= as7;
//         bs8 <= bs7;
//         cs8 <= cs7;
//         macs8 <= macs7;
//         as9 <= as8;
//         bs9 <= bs8;
//         cs9 <= cs8;
//         macs9 <= macs8;
//         as10 <= as9;
//         bs10 <= bs9;
//         cs10 <= cs9;
//         macs10 <= macs9;
//     endrule

//     rule rl_finish;
//        Bit#(32) mac_result = mac.get();
//       // if(count%12==0) 
//        // begin
//             if ((mac_result!=macs1)) 
//             begin
//                 //if(count>=7)
//                     failed_cases <= failed_cases + 1;
//                // $display("%d --Expected O/P --- %b, Actual O/P-- %b",count,pack(as10*bs10+cs10), mac_result);
//             end
//             if(count>=7)
//                 $display("%d A: %b  B: %b  C:%b \n--Expected O/P --- %b, Actual O/P-- %b",count,pack(as10),pack(bs10),pack(cs10),pack(macs1), mac_result);
//        // end
//         if(count==1060)
//             begin
//             $display("Failed for %d cases", failed_cases);
//             $finish(0);
//             end

//     endrule
//  endmodule



// (*always_ready*)
//   interface Ifc_inp;
//     method Action put_r( Bit#(1) read);
//     method Bit#(8) get_a;   
//     method Bit#(8) get_b;
//     method Bit#(32) get_c;
//     method Bit#(32) get_mac;
//   endinterface

//   import "BVI" file_read = 
//   module mk_inp_read ( Ifc_inp ) ;

//     method out_a get_a;
//     method out_b get_b;
//     method out_c get_c;
//     method out_mac get_mac;
//     method put_r(read) enable(EN);

//     default_clock clk(clk, (*unused*) CLK_GATE);
//     //default_reset rst(rst);
//     schedule (put_r) CF (get_a);
//     schedule (put_r) CF (get_b);
//     schedule (put_r) CF (get_c);
//     schedule (put_r) CF (get_mac);

//   endmodule

    module mk_int8_mac(Ifc_int8);
        Reg#(Bit#(8))       rg_a    <-  mkReg(?);
        Reg#(Bit#(8))       rg_b    <-  mkReg(?);
        Reg#(Bit#(32))      rg_c    <-  mkReg(?);
        Reg#(Bit#(32))      out     <-  mkReg(?);
        Reg#(Int#(32))      cyc     <-  mkReg(-1);
        Reg#(Bit#(16))      p1      <-  mkReg(?);

        Ifc_signedMul8 obj_mul <- mk_signed_mul8;

        rule r1(cyc<6 && cyc>0);
            cyc <= cyc+1;
        endrule

        rule r2(cyc==6);
            Bit#(16) prod = obj_mul.get();
            p1 <= prod;
            cyc <= cyc+1;
        endrule

        rule r3(cyc==7);
            Bit#(5) s1,s2,s3,s4,s5,s6,s7,s8;
            s1 = func_CLA(p1[3:0],rg_c[3:0],1'b0);
            s2 = func_CLA(p1[7:4],rg_c[7:4],s1[4]);
            s3 = func_CLA(p1[11:8],rg_c[11:8],s2[4]);
            s4 = func_CLA(p1[15:12],rg_c[15:12],s3[4]);
            s5 = func_CLA({p1[15],p1[15],p1[15],p1[15]},rg_c[19:16],s4[4]);
            s6 = func_CLA({p1[15],p1[15],p1[15],p1[15]},rg_c[23:20],s5[4]);
            s7 = func_CLA({p1[15],p1[15],p1[15],p1[15]},rg_c[27:24],s6[4]);
            s8 = func_CLA({p1[15],p1[15],p1[15],p1[15]},rg_c[31:28],s7[4]);

            out <= {s8[3:0],s7[3:0],s6[3:0],s5[3:0],s4[3:0],s3[3:0],s2[3:0],s1[3:0]};
            
            cyc <= 0;
        endrule

        rule disp;
            $display("output is :%b",out);
        endrule
        

        method Action       put(Bit#(8) a, Bit#(8) b, Bit#(32) c);
            rg_a <= a;
            rg_b <= b;
            rg_c <= c;
            cyc  <= 1;
            obj_mul.put_inp(a,b);
        endmethod


        method Bit#(32)     get();
            if(cyc==0)
                    return out;
            else
                    return 32'd0;
                    
        endmethod
    endmodule


    interface Ifc_signedMul8;
        method Action put_inp(Bit#(8) a, Bit#(8) b);
        method Bit#(16)     get();
    endinterface

    module mk_signed_mul8(Ifc_signedMul8) provisos(Bitwise#(Bit#(8)));

        Reg#(Bit#(8)) x <- mkReg(?);
        Reg#(Bit#(8)) y <- mkReg(?);
        Reg#(Bit#(16)) z <- mkReg(?);
       
        //REGISTERS FOR STORING STAGE 1 RESULTS
        Reg#(Bit#(1)) pp00 <- mkReg(0); 
        Reg#(Bit#(1)) pp01 <- mkReg(0);
        Reg#(Bit#(1)) pp10 <- mkReg(0);
        Reg#(Bit#(1)) pp07 <- mkReg(0);
        Reg#(Bit#(1)) pp16 <- mkReg(0);
        Reg#(Bit#(1)) pp21 <- mkReg(0);
        Reg#(Bit#(1)) pp30 <- mkReg(0);
        Reg#(Bit#(1)) pp35 <- mkReg(0);
        Reg#(Bit#(1)) pp41 <- mkReg(0);
        Reg#(Bit#(1)) pp50 <- mkReg(0);
        Reg#(Bit#(1)) pp57 <- mkReg(0);
        Reg#(Bit#(1)) pp77 <- mkReg(0);


        Reg#(Bit#(5)) s11 <- mkReg(0); 
        Reg#(Bit#(5)) s12 <- mkReg(0);
        Reg#(Bit#(5)) s13 <- mkReg(0);
        Reg#(Bit#(5)) s14 <- mkReg(0);
        Reg#(Bit#(5)) s15 <- mkReg(0);
        Reg#(Bit#(5)) s16 <- mkReg(0);
           
        //REGISTERS FOR STORING STAGE 2 RESULTS 
        Reg#(Bit#(1)) pp00_s2 <- mkReg(0); 
        Reg#(Bit#(1)) pp10_s2 <- mkReg(0);
        Reg#(Bit#(1)) pp01_s2 <- mkReg(0);
        Reg#(Bit#(1)) pp35_s2 <- mkReg(0);
        Reg#(Bit#(1)) pp57_s2 <- mkReg(0);
        Reg#(Bit#(1)) pp77_s2 <- mkReg(0);

        Reg#(Bit#(5)) s21 <- mkReg(0); 
        Reg#(Bit#(5)) s22 <- mkReg(0); 
        Reg#(Bit#(5)) s23 <- mkReg(0);   

        Reg#(Bit#(5)) s15_s2 <- mkReg(0); 
        Reg#(Bit#(5)) s11_s2 <- mkReg(0); 
        Reg#(Bit#(5)) s16_s2 <- mkReg(0);   

        //REGISTER FOR STORING STAGE 3 RESULTS
        Reg#(Bit#(2)) s31 <- mkReg(0);
        Reg#(Bit#(2)) s32 <- mkReg(0); 
        Reg#(Bit#(2)) s33 <- mkReg(0); 
        Reg#(Bit#(2)) s34 <- mkReg(0); 
        Reg#(Bit#(2)) s35 <- mkReg(0); 
        Reg#(Bit#(2)) s36 <- mkReg(0); 

        Reg#(Bit#(1)) pp00_s3         <-       mkReg(0);
        Reg#(Bit#(1)) pp01_s3         <-       mkReg(0);
        Reg#(Bit#(1)) pp10_s3         <-       mkReg(0);
        Reg#(Bit#(1)) pp77_s3         <-       mkReg(0);
        Reg#(Bit#(5)) s11_s3          <-       mkReg(0);
        Reg#(Bit#(5)) s16_s3          <-       mkReg(0);
        Reg#(Bit#(5)) s21_s3          <-       mkReg(0);
        Reg#(Bit#(5)) s22_s3          <-       mkReg(0);
        Reg#(Bit#(5)) s23_s3          <-       mkReg(0);

        //REGISTERS FOR STORING STAGE 4 RESULTS   
        Reg#(Bit#(5)) s41           <- mkReg(0); 
        Reg#(Bit#(5)) s42           <- mkReg(0);
        Reg#(Bit#(5)) s43           <- mkReg(0);
        Reg#(Bit#(5)) s44           <- mkReg(0);      
        Reg#(Bit#(1)) pp00_s4         <-       mkReg(0);

        rule stage1;
            Bit#(8) pp0,pp1,pp2,pp3,pp4,pp5,pp6,pp7;
            //PARTIAL PRODUCTS CALCULATION:
            pp0             =       {(~((x[7])&(y[0]))),((x[6:0])&(signExtend(y[0])))};
            pp1             =       {(~((x[7])&(y[1]))),((x[6:0])&(signExtend(y[1])))};
            pp2             =       {(~((x[7])&(y[2]))),((x[6:0])&(signExtend(y[2])))};
            pp3             =       {(~((x[7])&(y[3]))),((x[6:0])&(signExtend(y[3])))};
            pp4             =       {(~((x[7])&(y[4]))),((x[6:0])&(signExtend(y[4])))};
            pp5             =       {(~((x[7])&(y[5]))),((x[6:0])&(signExtend(y[5])))};
            pp6             =       {(~((x[7])&(y[6]))),((x[6:0])&(signExtend(y[6])))};
            pp7             =       {((x[7])&(y[7])),(~((x[6:0])&(signExtend(y[7]))))};

            //STAGE 1 REDUCTION:
            s11             <=       func_CLA(pp0[5:2],pp1[4:1],pp2[0]);
            s12             <=       func_CLA(pp2[5:2],pp3[4:1],pp4[0]);
            s13             <=       func_CLA(pp4[5:2],pp5[4:1],pp6[0]);
            s14             <=       func_CLA({pp6[3:1],pp0[6]},{pp7[2:0],pp1[5]},1'b0);
            s15             <=       func_CLA({pp4[7],pp3[7],pp2[7],pp1[7]},{pp5[6],pp4[6],pp3[6],pp2[6]},1'b1);
            s16             <=       func_CLA(pp6[7:4],pp7[6:3],pp5[5]);

            pp00            <=       pp0[0];
            pp01            <=       pp0[1];
            pp10            <=       pp1[0];
            pp07            <=       pp0[7];
            pp16            <=       pp1[6];
            pp21            <=       pp2[1];
            pp30            <=       pp3[0];
            pp35            <=       pp3[5];
            pp41            <=       pp4[1];
            pp50            <=       pp5[0];
            pp57            <=       pp5[7];
            pp77            <=       pp7[7];
        endrule

        rule stage2;
            //STAGE 2 REDUCTION:
            s21             <=       func_CLA(s11[4:1],{s12[2:0],pp21},pp30);
            s22             <=       func_CLA({s13[2:0],pp41},{s14[2:0],pp50},1'b0);
            s23             <=       func_CLA({s13[4:3],s15[0],pp07},{s14[4:3],s12[4:3]},pp16);

            pp00_s2         <=       pp00;
            pp01_s2         <=       pp01;
            pp10_s2         <=       pp10;
            pp35_s2         <=       pp35;
            pp57_s2         <=       pp57;
            pp77_s2         <=       pp77;
            s15_s2          <=       s15;
            s11_s2          <=       s11;
            s16_s2          <=       s16;

        endrule

        rule stage3;

            Bit#(2) temp1,temp2,temp3,temp4,temp5,temp6;
            //STAGE 3 REDUCTION:
            temp1           =       func_HA(s21[4],s22[2]);
            temp2           =       func_FA(pp35_s2,s22[3],s23[1]);
            temp3           =       func_FA(s15_s2[1],s22[4],s23[2]);
            temp4           =       func_FA(s15_s2[2],s16_s2[0],s23[3]);
            temp5           =       func_FA(s15_s2[3],s16_s2[1],s23[4]);
            temp6           =       func_FA(s15_s2[4],s16_s2[2],pp57_s2);

            s31             <=      {temp1[0],temp1[1]};
            s32             <=      {temp2[0],temp2[1]};
            s33             <=      {temp3[0],temp3[1]};
            s34             <=      {temp4[0],temp4[1]};
            s35             <=      {temp5[0],temp5[1]};
            s36             <=      {temp6[0],temp6[1]};

            pp00_s3         <=       pp00_s2;
            pp01_s3         <=       pp01_s2;
            pp10_s3         <=       pp10_s2;
            pp77_s3         <=       pp77_s2;
            s11_s3          <=       s11_s2;
            s16_s3          <=       s16_s2;
            s21_s3          <=       s21;
            s22_s3          <=       s22;
            s23_s3          <=       s23;
        endrule

        rule stage4;
            //VECTOR MERGE STAGE:
            s41             <=       func_CLA({s21_s3[1:0],s11_s3[0],pp01_s3},{3'b0,pp10_s3},1'b0);
            s42             <=       func_CLA({s32[0],s31[0],s21_s3[3:2]},{s31[1],s23_s3[0],s22_s3[1:0]},s41[4]);
            s43             <=       func_CLA({s36[0],s35[0],s34[0],s33[0]},{s35[1],s34[1],s33[1],s32[1]},s42[4]);
            s44             <=       func_CLA({1'b0,1'b1,pp77_s3,s16[3]},{2'b0,s16_s3[4],s36[1]},s43[4]);

            pp00_s4         <=       pp00_s3;

        endrule

        rule res1;
             Bit#(16) z_out = {s44[2],s44[1],s44[0],s43[3],s43[2],s43[1],s43[0],s42[3],s42[2],s42[1],s42[0],s41[3],s41[2],s41[1],s41[0],pp00_s4};
             z <= z_out;
        endrule


        method Action put_inp(Bit#(8) a, Bit#(8) b);
            x <= a;
            y <= b;
        endmethod

        method Bit#(16)     get();
            return z;
        endmethod

    endmodule



    //1. 4-bit Carry Lookahead Adder
    function Bit#(5) func_CLA(Bit#(4) rg_a, Bit#(4) rg_b, bit cin);
        Bit#(4)             g,p,sum,carrrg_b;
        bit                 cout;
        g               =   rg_a&rg_b;
        p               =   rg_a^rg_b;
        carrrg_b[0]     =   cin;
        carrrg_b[1]     =   g[0] | p[0]&cin;
        carrrg_b[2]     =   g[1] | p[1]&g[0] | p[1]&p[0]&cin;
        carrrg_b[3]     =   g[2] | p[2]&g[1] | p[2]&p[1]&g[0] | p[2]&p[1]&p[0]&cin;
        cout            =   g[3] | p[3]&g[2] | p[3]&p[2]&g[1] | p[3]&p[2]&p[1]&g[0] | p[3]&p[2]&p[1]&p[0]&cin; 
        sum             =   p ^ carrrg_b;
        return    {cout, sum};
    endfunction

    //2. Half Adder
    function Bit#(2) func_HA(bit a, bit b);
        Bit#(2) sum;
        sum[1]          =   a^b;
        sum[0]          =   a&b;
        return sum;
    endfunction

    //3. Full Adder
    function Bit#(2) func_FA(bit a, bit b, bit cin);
        Bit#(2) sum;
        sum[1]          =   a^b^cin;
        sum[0]          =   (a&b) | (a^b)&cin;
        return sum;
    endfunction
endpackage